module write_back_phase (
    input logic writeback
    
);
    
endmodule