module write_back_phase (
    
);
    
endmodule